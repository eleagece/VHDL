library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-------------------------------------------------------------------------------------------------------
-- Entity memoria
-------------------------------------------------------------------------------------------------------
entity memoria is
	port ( clk: in std_logic;
			 reset: in std_logic; -- borra la memoria
			 en: in std_logic; -- enable
			 l: in std_logic; -- leer 1
			 e: in std_logic; -- escribir 1
			 dataIn: in std_logic_vector(8 downto 0); -- valor RGB para meter
			 dataOut: out std_logic_vector(8 downto 0); -- valor RGB para sacar
			 dir: in std_logic_vector(6 downto 0) ); -- selecciona una de las 128 posiciones para leer o escribir
end memoria;

-------------------------------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------------------------------
architecture Behavioral of memoria is

--> Types, signals
type tipo is array(0 to 127) of std_logic_vector(8 downto 0);
signal datos: tipo:=("111000000","111000000","110000000","110000000",
							"101000000","101000000","100000000","100000000", 
							"011000000","011000000","010000000","010000000", -- linea 1
							"001000000","001000000","001000000","001000000", -- 0-15
							
							"111000000","111111111","110000000","111111111",
							"101000000","111111111","100000000","111111111",
							"011000000","111111111","111111111","010000000", -- linea 2
							"001000000","111111111","001000000","001000000", -- 16-31
							
							"111000000","111111111","110000000","111111111",
							"101000000","111111111","100000000","111111111", 
							"011000000","111111111","010000000","111111111", -- linea 3
							"001000000","111111111","001000000","001000000", -- 32-47
							
							"111000000","111111111","110000000","111111111",
							"101000000","111111111","111111111","111111111",
							"011000000","111111111","010000000","111111111", -- linea 4
							"001000000","111111111","001000000","001000000", -- 48-63
							
							"111000000","111111111","110000000","111111111",
							"101000000","111111111","111111111","111111111",
							"011000000","111111111","010000000","111111111", -- linea 5
							"001000000","111111111","001000000","001000000", -- 64-79
							
							"111000000","111111111","110000000","111111111",
							"101000000","111111111","100000000","111111111",
							"011000000","111111111","010000000","111111111", -- linea 6
							"001000000","111111111","001000000","001000000", -- 80-95
							
							"111000000","111000000","111111111","110000000", 
							"101000000","111111111","100000000","111111111",
							"011000000","111111111","111111111","010000000", -- linea 7
							"001000000","111111111","111111111","001000000", -- 96-111
							
							"111000000","111000000","110000000","110000000",
							"101000000","101000000","100000000","100000000", 
							"011000000","011000000","010000000","010000000", -- linea 8
							"001000000","001000000","001000000","001000000"); -- 112-127               
							
--> Begin architecture
begin

-->> Process
-->>> Proceso de reseteo, lectura y escritura en memoria
process(l,e,en,clk)
begin
	if (en='1') then
		if (clk'event and clk='1') then
			if (e='1' and l='0') then
				datos(conv_integer(dir))<=dataIn;
			elsif (e='0' and l='1') then
				dataOut<=datos(conv_integer(dir));
			else
				dataOut<="111000000";
			end if;
		end if;
	else
		dataOut<="111000000";
	end if;
end process;

end Behavioral;
