library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-------------------------------------------------------------------------------------------------------
-- Entity vgacore
-------------------------------------------------------------------------------------------------------
entity vgacore is
	port ( reset: in std_logic; -- reset
		    clock: in std_logic; -- reloj de la FPGA a 100 Mhz
			 weRX: in std_logic; -- llega dato nuevo
			 recibir: in std_logic; -- permite recibir un mensaje
			 doutRX: in std_logic_vector(5 downto 0); -- dato actualmente le�do de la memoria
		    hsyncb: inout std_logic; -- horizontal (line) sync
		    vsyncb: out std_logic;	-- vertical (frame) sync
		    rgb: out std_logic_vector(8 downto 0) ); -- red, green, blue colores
end vgacore;

-------------------------------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------------------------------
architecture vgacore_arch of vgacore is

-- Components -----------------------------------------------------------------------------------------

-- Types, constants, signals --------------------------------------------------------------------------
-->> vgacore pantalla
signal hcnt: std_logic_vector(8 downto 0); -- horizontal pixel counter
signal vcnt: std_logic_vector(9 downto 0); -- vertical line counter

-->> vgacore reloj pantalla
signal contadorClk: std_logic_vector(1 downto 0); -- contador para dividir la frecuencia del contador interno
signal clk: std_logic; -- reloj de la pantalla (12,5 Mhz)

-->> m�quina de estados
type TEstado is (ESPERA,R0,R1,R2); 
signal estado,nestado:TEstado;

-->> cuenta interno
signal cuenta: std_logic_vector(6 downto 0); -- �ndice por el que vamos del mensaje
signal ncuenta: std_logic_vector(6 downto 0);
signal glscene: std_logic;

-->> ram que guarda los valores del mensaje, los cuales act�an de �ndice de arrayLetrasDesp para hallar el desplazamiento
type arrayBaseLetra is array(0 to 127) of std_logic_vector(5 downto 0);
signal baseLetra: arrayBaseLetra:=(others=>"000000");
-- (0=>"000000", 1=>"000001", 2=>"000010", 3=>"000011", 4=>"000100", 
--  5=>"000101", 6=>"000110", 7=>"000111", 8=>"001000", 9=>"001001", 
--  10=>"001010", 11=>"001011", 12=>"001100", 13=>"001101", 14=>"001110", 
--  15=>"001111", 16=>"010000", 17=>"010001", 18=>"010010", 19=>"010011",
--  20=>"010100", 21=>"010101", 22=>"010110", 23=>"010111", 24=>"011000",
--  25=>"011001", 26=>"011010", 27=>"011011", 28=>"011100", 29=>"011101", 
--  30=>"011110", 31=>"011111", 32=>"100000", 33=>"100001", 34=>"100010",
--  35=>"100011", 36=>"100100", others=>"000000");

-->> roms de sprites de letras
type arraySpriteLetras is array(0 to 15) of std_logic_vector(7 downto 0);
signal filaSpriteLetras: arraySpriteLetras; -- array que guarda 0, 8, 8+8, 8+8+8... para sacar la posici�n en memoria de cada fila de la letra
type arrayLetrasDesp is array(0 to 36) of std_logic_vector(12 downto 0); 
signal posicionLetrasDesp: arrayLetrasDesp; -- array que guarda 0, 128, 128+128... para sacar la posici�n en memoria de cada letra
type spriteLetras is array(0 to 4735) of std_logic; -- p�xeles de las letras del mensaje
signal letras: spriteLetras:=
	-- 0
	('0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','1','0','1','0','0','0','1',
	 '0','1','0','1','0','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	-- 1
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','1','1','0','0',
	 '0','0','0','0','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','1','1','1','1','1',
	 '0','0','0','1','1','1','1','1',
	-- 2
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','0','1','1','1','1','0',
	 '0','0','0','1','1','1','1','0',
	 '0','0','1','0','0','0','0','0',
	 '0','0','1','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	-- 3
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- 4
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	-- 5
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	-- 6
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	-- 7
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	-- 8
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- 9
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- A
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- B
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	-- C
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	-- D
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	-- E
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	-- F
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	-- G
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','1','1','1',
	 '0','1','0','0','0','1','1','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- H
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- I
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','1','1','1','0','0',
	 '0','0','0','1','1','1','0','0',
	-- J
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','1','1','1',
	 '0','0','0','0','0','1','1','1',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','1','0','0','0','0','1','0',
	 '0','1','0','0','0','0','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- K
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','1','1',
	 '0','1','0','0','0','0','1','1',
	 '0','1','0','0','0','1','0','0',
	 '0','1','0','0','0','1','0','0',
	 '0','1','0','0','1','0','0','0',
	 '0','1','0','0','1','0','0','0',
	 '0','1','1','1','0','0','0','0',
	 '0','1','1','1','0','0','0','0',
	 '0','1','0','0','1','0','0','0',
	 '0','1','0','0','1','0','0','0',
	 '0','1','0','0','0','1','0','0',
	 '0','1','0','0','0','1','0','0',
	 '0','1','0','0','0','0','1','1',
	 '0','1','0','0','0','0','1','1',
	-- L
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	-- M
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','0','0','0','1','1',
	 '0','1','1','0','0','0','1','1',
	 '0','1','1','1','0','1','1','1',
	 '0','1','1','1','0','1','1','1',
	 '0','1','0','1','0','1','0','1',
	 '0','1','0','1','0','1','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- N
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','0','0','0','0','1',
	 '0','1','1','0','0','0','0','1',
	 '0','1','0','1','0','0','0','1',
	 '0','1','0','1','0','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','1','0','0','0','0','1','1',
	 '0','1','0','0','0','0','1','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- O
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- P
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	-- Q
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','1','0','0','0','1','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- R
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- S
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','1',
	 '0','0','1','1','1','1','1','1',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','0','0','0','0','0','0','1',
	 '0','1','1','1','1','1','1','0',
	 '0','1','1','1','1','1','1','0',
	-- T
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	-- U
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','1','1','1','1','0',
	 '0','0','1','1','1','1','1','0',
	-- V
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','1','0',
	 '0','1','0','0','0','0','1','0',
	 '0','0','1','0','0','1','0','0',
	 '0','0','1','0','0','1','0','0',
	 '0','0','0','1','1','0','0','0',
	 '0','0','0','1','1','0','0','0',
	-- W
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','0','1','0','0','1',
	 '0','1','0','1','0','1','0','1',
	 '0','1','0','1','0','1','0','1',
	 '0','1','1','0','0','0','1','1',
	 '0','1','1','0','0','0','1','1',
	-- X
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	-- Y
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','0','0','0','0','0','1',
	 '0','1','0','0','0','0','0','1',
	 '0','0','1','0','0','0','1','0',
	 '0','0','1','0','0','0','1','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','0','1','0','1','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	-- Z
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','0','1','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','0','1','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','0','1','0','0','0',
	 '0','0','0','1','0','0','0','0',
	 '0','0','0','1','0','0','0','0',
	 '0','0','1','0','0','0','0','0',
	 '0','0','1','0','0','0','0','0',
	 '0','1','1','1','1','1','1','1',
	 '0','1','1','1','1','1','1','1',
	-- ESPACIO
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0',
	 '0','0','0','0','0','0','0','0');

--type spriteMorse is array(0 to 21887) of std_logic; -- p�xeles de las letras en morse del mensaje
--type arraySpriteMorse is array(0 to 575) of std_logic_vector(CALCULAR TAMA�O downto 0);
--signal filaSpriteMorse: arraySpriteMorse; -- array que guarda 0, 38, 38+38, 38+38+38... para sacar la posici�n en memoria de cada fila
--signal morse: spriteMorse:=
--     (PONER LA CODIFICACI�N DE LAS LETRAS EN MORSE);
	  
-------------------------------------------------------------------------------------------------------
-- Begin architecture
-------------------------------------------------------------------------------------------------------
begin

-- Combinacional --------------------------------------------------------------------------------------
-->> empty

-- Generates ------------------------------------------------------------------------------------------
-->> generate que indica la fila por la que se va pintando la letra
filaSpriteLetras(0)<=(others=>'0');
gen1: for i in 1 to 15 generate
	filaSpriteLetras(i)<=filaSpriteLetras(i-1)+"00001000";
end generate gen1;

posicionLetrasDesp(0)<=(others=>'0');
gen2: for i in 1 to 36 generate
	posicionLetrasDesp(i)<=posicionLetrasDesp(i-1)+"10000000";
end generate gen2;

-- Component port maps --------------------------------------------------------------------------------
-->> empty

-- Process --------------------------------------------------------------------------------------------
-->> proceso A: aumenta hcnt con cada ciclo de reloj desde 0 a 380 y lo vuelve a 0.
A: process(clk,reset)
begin
	-- reset asynchronously clears pixel counter
	if reset='1' then
		hcnt <= "000000000";
	-- horiz. pixel counter increments on rising edge of dot clk
	elsif (clk'event and clk='1') then
		-- horiz. pixel counter rolls-over after 381 pixels
		if hcnt<380 then
			hcnt <= hcnt + 1;
		else
			hcnt <= "000000000";
		end if;
	end if;
end process;

-->> proceso B: aumenta vcnt con cada ciclo de hsyncb desde 0 a 527 y lo vuelve a 0.
B: process(hsyncb,reset)
begin
	-- reset asynchronously clears line counter
	if reset='1' then
		vcnt <= "0000000000";
	-- vert. line counter increments after every horiz. line
	elsif (hsyncb'event and hsyncb='1') then
		-- vert. line counter rolls-over after 528 lines
		if vcnt<527 then
			vcnt <= vcnt + 1;
		else
			vcnt <= "0000000000";
		end if;
	end if;
end process;

-->> proceso C
C: process(clk,reset)
begin
	-- reset asynchronously sets horizontal sync to inactive
	if reset='1' then
		hsyncb <= '1';
	-- horizontal sync is recomputed on the rising edge of every dot clk
	elsif (clk'event and clk='1') then
		-- horiz. sync is low in this interval to signal start of a new line
		if (hcnt>=291 and hcnt<337) then
			hsyncb <= '0';
		else
			hsyncb <= '1';
		end if;
	end if;
end process;

-->> proceso D
D: process(hsyncb,reset)
begin
	-- reset asynchronously sets vertical sync to inactive
	if reset='1' then
		vsyncb <= '1';
	-- vertical sync is recomputed at the end of every line of pixels
	elsif (hsyncb'event and hsyncb='1') then
		-- vert. sync is low in this interval to signal start of a new frame
		if (vcnt>=490 and vcnt<492) then
			vsyncb <= '0';
		else
			vsyncb <= '1';
		end if;
	end if;
end process;

-->> proceso que consigue el reloj de 12,5 Mhz al que funciona la pantalla
process (reset,clock,contadorClk)
begin
	if (reset='1') then
		contadorClk<="00";
		clk<='0';
	elsif clock'event and clock='1' then
		if (contadorClk="11") then
			clk<=not clk;
			contadorClk<="00";
		else
			contadorClk<=contadorClk+1;
		end if;
	end if;
end process;

-->> Proceso de cambio de estado
process(clk,reset)
begin
	if reset='1' then 
		estado<=ESPERA;
		cuenta<=(others=>'0');
	elsif clk'event and clk='1' then
		cuenta<=ncuenta;
		estado<=nestado;
	end if;
end process;

-->> Proceso de gu�a de cambio de estado
process (estado,recibir,weRX,clk,cuenta)
begin
	nestado<=estado;
	ncuenta<=cuenta;
	glscene<='0';
	case estado is
	 -- estado ESPERA
		when ESPERA=>
			if (recibir='1') then
				nestado<=R0;
			end if;
	 -- estados de recibir
		when R0=>
			if recibir='0' then
				nestado<=ESPERA;
				ncuenta<=(others=>'0');
			elsif (weRX='1') then
				nestado<=R1;
				ncuenta<=cuenta+1;
			end if;
		when R1=>
			glscene<='1';
			nestado<=R2;
		when R2=>
			if (weRX='0') then
				nestado<=R0;
			end if;
	end case;			
end process;

process(glscene,clk,reset)
	begin
		if reset='1' then
				baseLetra(0)<="100100";
		elsif (clk'event and clk='1') then
			if glscene='1' then
				baseLetra(conv_integer(cuenta))<=doutRX;
			else
				baseLetra(conv_integer(cuenta))<=baseLetra(conv_integer(cuenta));
			end if;
		end if; 
	end process;

-->> Proceso de dibujado
process(vcnt,hcnt)
begin
	rgb<=(others=>'0');
	-- marco de recibir
	if ((vcnt=16) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=16
		((vcnt=45) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=45
		((vcnt>=16 and vcnt<46) and (hcnt=254)) xor -- vertical (16 a 45) en hcnt=254
		((vcnt>=16 and vcnt<46) and (hcnt=283)) then -- vertical (16 a 45) en hcnt=283;
		if (modo='recibir')
			rgb<="000111000";
		else
			rgb<="111111111";
		end if
	-- letra de recibir
	elsif (hcnt>=266 and hcnt<=273 and vcnt>=22 and vcnt<=37) then
		if (letras(conv_integer( filaSpriteLetras(conv_integer(vcnt-22)) + (hcnt-266) + 3456))='1')
			if (modo='recibir')
				rgb<="000111000";
			else
				rgb<="111111111";
			end if;
		else
			rgb<=(others=>'0');
		end if;
	-- marco de escribir
	elsif ((vcnt=57) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=57
		((vcnt=86) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=86
		((vcnt>=57 and vcnt<87) and (hcnt=254)) xor -- vertical (57 a 86) en hcnt=254
		((vcnt>=57 and vcnt<87) and (hcnt=283)) then -- vertical (57 a 86) en hcnt=283
		if (modo='escribir')
			rgb<="000111000";
		else
			rgb<="111111111";
		end if
	-- letra de escribir
	elsif (hcnt>=266 and hcnt<=273 and vcnt>=63 and vcnt<=78) then
		if (letras(conv_integer( filaSpriteLetras(conv_integer(vcnt-63)) + (hcnt-266) + 1792))='1')
			if (modo='escribir')
				rgb<="000111000";
			else
				rgb<="111111111";
			end if;
		else
			rgb<=(others=>'0');
		end if;
	-- marco de transmitir
	elsif ((vcnt=98) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=98
		((vcnt=127) and (hcnt>254 and hcnt<282)) xor -- horizontal (255 a 282) en vcnt=127
		((vcnt>=98 and vcnt<128) and (hcnt=254)) xor -- vertical (98 a 127) en hcnt=254
		((vcnt>=98 and vcnt<128) and (hcnt=283)) then -- vertical (98 a 127) en hcnt=283
		if (modo='transmitir')
			rgb<="000111000";
		else
			rgb<="111111111";
		end if
	-- letra de transmitir
	elsif (hcnt>=266 and hcnt<=273 and vcnt>=104 and vcnt<=119) then
		if (letras(conv_integer( filaSpriteLetras(conv_integer(vcnt-104)) + (hcnt-266) + 3712))='1')
			if (modo='transmitir')
				rgb<="000111000";
			else
				rgb<="111111111";
			end if;
		else
			rgb<=(others=>'0');
		end if;
	-- marco del mensaje
	elsif ((vcnt=0) and (hcnt>0 and hcnt<289)) xor -- horizontal (1 a 288) en vcnt=0
		((vcnt=144) and (hcnt>0 and hcnt<289)) xor -- horizontal (1 a 288) en vcnt=144
		((vcnt>=0 and vcnt<145) and (hcnt=0)) xor -- vertical (0 a 144) en hcnt=0
		((vcnt>=0 and vcnt<145) and (hcnt=289)) then -- vertical (0 a 144) en hcnt=289
		rgb<=(others=>'1');
	-- mensaje
	elsif (hcnt>7 and hcnt<248) then
		if (vcnt>15 and vcnt<32) then
			if (letras(conv_integer(posicionLetrasDesp(conv_integer(baseLetra(conv_integer(hcnt(7 downto 3))-1))) + filaSpriteLetras(conv_integer(vcnt(3 downto 0))) + hcnt(2 downto 0)))='1') then
					--and (hcnt(7 downto 3))<=cuenta) then
				rgb<=(others=>'1');
			end if;
		elsif (vcnt>47 and vcnt<64) then
			if (letras(conv_integer(posicionLetrasDesp(conv_integer(baseLetra(conv_integer(hcnt(7 downto 3))+29))) + filaSpriteLetras(conv_integer(vcnt(3 downto 0))) + hcnt(2 downto 0)))='1') then
					--and ((hcnt(7 downto 3))+32)<=cuenta) then
				rgb<=(others=>'1');
			end if;
		elsif (vcnt>79 and vcnt<96) then
			if (letras(conv_integer(posicionLetrasDesp(conv_integer(baseLetra(conv_integer(hcnt(7 downto 3))+59))) + filaSpriteLetras(conv_integer(vcnt(3 downto 0))) + hcnt(2 downto 0)))='1') then
					--and ((hcnt(7 downto 3))+64)<=cuenta) then
				rgb<=(others=>'1');
			end if;
		elsif (vcnt>111 and vcnt<128) then
			if (letras(conv_integer(posicionLetrasDesp(conv_integer(baseLetra(conv_integer(hcnt(7 downto 3))+89))) + filaSpriteLetras(conv_integer(vcnt(3 downto 0))) + hcnt(2 downto 0)))='1') then
					--and ((hcnt(7 downto 3))+96)<=cuenta) then
				rgb<=(others=>'1');
			end if;
		end if;
	end if;
end process;

end vgacore_arch;

